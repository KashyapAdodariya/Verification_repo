

// Revision: 1
//-------------------------------------------------------------------------------

package pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

`include "cfg.sv"
`include "report_catcher.sv"
//`include "report_server.sv"
`include "sequence_item.sv"
`include "coverage.sv"
`include "callback_comp.sv"
`include "callback_seq.sv"
`include "reg_block.sv"
`include "ral_adepter.sv"
`include "env_cfg.sv"
`include "agent_cfg.sv"
`include "slave_mem.sv"
`include "sequencer.sv"
`include "slave_seqr.sv"
`include "sequence.sv"
`include "slave_seq.sv"
`include "virtual_seqr.sv"
`include "scoreboard.sv"
`include "driver.sv"
`include "slave_drv.sv"
`include "monitor.sv"
`include "slave_mon.sv"
`include "agent.sv"
`include "slave_agt.sv"
`include "ral_env.sv"
`include "env.sv"
`include "virtual_seq.sv"
`include "test.sv"
  
endpackage:pkg


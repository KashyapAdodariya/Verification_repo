Example for UVM callback in uvm_sequence
Run Options: +UVM_TESTNAME=base_test
Run Options: +UVM_TESTNAME=err_test
`include "seq_item.sv"
`include "all_reg_pkt.sv"
`include "ral_adapter.sv"
`include "sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "ral_env.sv"
`include "sys_env.sv"


//Used case of callback add method with two callback class
//if used `uvm_do_callbacks(...); then no matter which one excute first
/*package i2s_pkg;
 
  import uvm_pkg::*;
  `include "uvm_macros.svh"

endpackage:i2s_pkg
*/
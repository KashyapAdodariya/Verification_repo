

`define print(MSG) `uvm_info("DEMO-V0.2", MSG, UVM_LOW)
interface i2s_interface (input bit clk);
  logic a;
  //$display("i2s_interface run");
endinterface




package sv_pkg;

	`include "transaction_item.sv"
	`include "monitor.sv"
	`include "scb.sv"
	`include "scb_subscriber.sv"
	`include "scb_wrapper.sv"
	`include "env.sv"
	`include "test.sv"

endpackage: sv_pkg
interface intf_h(input bit clock);
  logic [7:0]addr;
  logic [31:0]data;
endinterface: intf_h
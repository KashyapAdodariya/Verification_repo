`include "axi_m_config.sv"
`include "axi_m_tran.sv"
`include "axi_m_tran.svh"
`include "axi_intf.sv"
`include "axi_m_monitor.sv"
`include "axi_m_scoreboard.sv"
`include "axi_m_gen.sv"
`include "axi_m_driver.sv"
`include "axi_s_dri.sv"
`include "axi_m_agent.sv"
`include "axi_m_env.sv"
`include "axi_m_tb.sv"

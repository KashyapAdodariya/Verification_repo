

`define print(MSG) `uvm_info(get_type_name(), MSG, UVM_LOW)